LIBRARY IEEE;
USE IEEE.std_logic_1164.all;
USE IEEE.numeric_std.all;
USE IEEE.std_logic_signed.all;

ENTITY RAM_ADDRESS_RESOLVER IS
		PORT( 
		SIZE: IN std_logic;
		READ_FILTER: IN std_logic;
		ROWS_COUNTER: IN std_logic_vector(7 DOWNTO 0);
		COLS_COUNTER: IN std_logic_vector(7 DOWNTO 0);
		RAM_ADDRESS_VALUE: IN std_logic_vector(17 DOWNTO 0);
		Q: OUT std_logic_vector(17 DOWNTO 0)
		);
END RAM_ADDRESS_RESOLVER;


ARCHITECTURE RAR_ARCH OF RAM_ADDRESS_RESOLVER IS

SIGNAL ADDRESS_VALUE: std_logic_vector(17 downto 0);

BEGIN
	
	PROCESS (READ_FILTER, ROWS_COUNTER, COLS_COUNTER, RAM_ADDRESS_VALUE)
	BEGIN
		IF (ROWS_COUNTER = "00000000") THEN
			IF (READ_FILTER = '1') THEN
				ADDRESS_VALUE <= (OTHERS => '0');
			ELSIF (SIZE = '0') THEN
				ADDRESS_VALUE <= "000000000000001001" + ("0000000000" & COLS_COUNTER);
			ELSE
				ADDRESS_VALUE <= "000000000000011001" + ("0000000000" & COLS_COUNTER);
			END IF;
		ELSIF (READ_FILTER = '1') THEN
		  IF (SIZE = '1') THEN
			   ADDRESS_VALUE <= RAM_ADDRESS_VALUE + "000000000000000101";
			ELSE 
			   ADDRESS_VALUE <= RAM_ADDRESS_VALUE + "000000000000000011";
			END IF;
		ELSE 
			ADDRESS_VALUE <= RAM_ADDRESS_VALUE + "000000000100000000";
		END IF;
	END PROCESS;

	Q <= ADDRESS_VALUE;	

END RAR_ARCH;

